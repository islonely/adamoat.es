module main

import veb

pub struct Context {
	veb.Context
}
